`timescale 1ns/1ns
module testbench;
    reg RESET;
    reg RXD;
    wire TXD;
    wire PWM;    

    SOC uut (
        .RESET(RESET), 
        .RXD(RXD),
        .TXD(TXD),
        .PWM(PWM)
    );

    initial begin
        $dumpfile("test.vcd");
        $dumpvars(0, testbench);

        // Init
        RXD = 1;
        RESET = 0;

        // Reset Pulse
        #100 RESET = 1;
        #100 RESET = 0; 

        #1000000000;
        $finish;
    end
endmodule
